`timescale 1ns / 1ps

module DFF(
    output reg q,
    output reg qBar,
    input d,
    input clk,
    input resetBar
    );

wire tmp0;
wire tmp1;
wire tmp2;
wire tmp3;


    always @ (tmp3) begin
        None <= tmp3;
    end


    always @ (tmp2) begin
        None <= tmp2;
    end


    always @ (tmp1) begin
        None <= tmp1;
    end


    always @ (tmp0) begin
        None <= tmp0;
    end


    always @ (qBar) begin
        None <= qBar;
    end


    always @ (q) begin
        None <= q;
    end

endmodule
